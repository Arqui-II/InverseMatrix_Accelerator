// Nios2_accelerator.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module Nios2_accelerator (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

	wire         nios_ii_custom_instruction_master_readra;                                      // NIOS_II:D_ci_readra -> NIOS_II_custom_instruction_master_translator:ci_slave_readra
	wire   [4:0] nios_ii_custom_instruction_master_a;                                           // NIOS_II:D_ci_a -> NIOS_II_custom_instruction_master_translator:ci_slave_a
	wire   [4:0] nios_ii_custom_instruction_master_b;                                           // NIOS_II:D_ci_b -> NIOS_II_custom_instruction_master_translator:ci_slave_b
	wire   [4:0] nios_ii_custom_instruction_master_c;                                           // NIOS_II:D_ci_c -> NIOS_II_custom_instruction_master_translator:ci_slave_c
	wire         nios_ii_custom_instruction_master_readrb;                                      // NIOS_II:D_ci_readrb -> NIOS_II_custom_instruction_master_translator:ci_slave_readrb
	wire         nios_ii_custom_instruction_master_clk;                                         // NIOS_II:E_ci_multi_clock -> NIOS_II_custom_instruction_master_translator:ci_slave_multi_clk
	wire  [31:0] nios_ii_custom_instruction_master_ipending;                                    // NIOS_II:W_ci_ipending -> NIOS_II_custom_instruction_master_translator:ci_slave_ipending
	wire         nios_ii_custom_instruction_master_start;                                       // NIOS_II:E_ci_multi_start -> NIOS_II_custom_instruction_master_translator:ci_slave_multi_start
	wire         nios_ii_custom_instruction_master_reset_req;                                   // NIOS_II:E_ci_multi_reset_req -> NIOS_II_custom_instruction_master_translator:ci_slave_multi_reset_req
	wire         nios_ii_custom_instruction_master_done;                                        // NIOS_II_custom_instruction_master_translator:ci_slave_multi_done -> NIOS_II:E_ci_multi_done
	wire   [7:0] nios_ii_custom_instruction_master_n;                                           // NIOS_II:D_ci_n -> NIOS_II_custom_instruction_master_translator:ci_slave_n
	wire  [31:0] nios_ii_custom_instruction_master_result;                                      // NIOS_II_custom_instruction_master_translator:ci_slave_result -> NIOS_II:E_ci_result
	wire         nios_ii_custom_instruction_master_estatus;                                     // NIOS_II:W_ci_estatus -> NIOS_II_custom_instruction_master_translator:ci_slave_estatus
	wire         nios_ii_custom_instruction_master_clk_en;                                      // NIOS_II:E_ci_multi_clk_en -> NIOS_II_custom_instruction_master_translator:ci_slave_multi_clken
	wire  [31:0] nios_ii_custom_instruction_master_datab;                                       // NIOS_II:E_ci_datab -> NIOS_II_custom_instruction_master_translator:ci_slave_datab
	wire  [31:0] nios_ii_custom_instruction_master_dataa;                                       // NIOS_II:E_ci_dataa -> NIOS_II_custom_instruction_master_translator:ci_slave_dataa
	wire         nios_ii_custom_instruction_master_reset;                                       // NIOS_II:E_ci_multi_reset -> NIOS_II_custom_instruction_master_translator:ci_slave_multi_reset
	wire         nios_ii_custom_instruction_master_writerc;                                     // NIOS_II:D_ci_writerc -> NIOS_II_custom_instruction_master_translator:ci_slave_writerc
	wire  [31:0] nios_ii_custom_instruction_master_translator_comb_ci_master_result;            // NIOS_II_custom_instruction_master_comb_xconnect:ci_slave_result -> NIOS_II_custom_instruction_master_translator:comb_ci_master_result
	wire         nios_ii_custom_instruction_master_translator_comb_ci_master_readra;            // NIOS_II_custom_instruction_master_translator:comb_ci_master_readra -> NIOS_II_custom_instruction_master_comb_xconnect:ci_slave_readra
	wire   [4:0] nios_ii_custom_instruction_master_translator_comb_ci_master_a;                 // NIOS_II_custom_instruction_master_translator:comb_ci_master_a -> NIOS_II_custom_instruction_master_comb_xconnect:ci_slave_a
	wire   [4:0] nios_ii_custom_instruction_master_translator_comb_ci_master_b;                 // NIOS_II_custom_instruction_master_translator:comb_ci_master_b -> NIOS_II_custom_instruction_master_comb_xconnect:ci_slave_b
	wire         nios_ii_custom_instruction_master_translator_comb_ci_master_readrb;            // NIOS_II_custom_instruction_master_translator:comb_ci_master_readrb -> NIOS_II_custom_instruction_master_comb_xconnect:ci_slave_readrb
	wire   [4:0] nios_ii_custom_instruction_master_translator_comb_ci_master_c;                 // NIOS_II_custom_instruction_master_translator:comb_ci_master_c -> NIOS_II_custom_instruction_master_comb_xconnect:ci_slave_c
	wire         nios_ii_custom_instruction_master_translator_comb_ci_master_estatus;           // NIOS_II_custom_instruction_master_translator:comb_ci_master_estatus -> NIOS_II_custom_instruction_master_comb_xconnect:ci_slave_estatus
	wire  [31:0] nios_ii_custom_instruction_master_translator_comb_ci_master_ipending;          // NIOS_II_custom_instruction_master_translator:comb_ci_master_ipending -> NIOS_II_custom_instruction_master_comb_xconnect:ci_slave_ipending
	wire  [31:0] nios_ii_custom_instruction_master_translator_comb_ci_master_datab;             // NIOS_II_custom_instruction_master_translator:comb_ci_master_datab -> NIOS_II_custom_instruction_master_comb_xconnect:ci_slave_datab
	wire  [31:0] nios_ii_custom_instruction_master_translator_comb_ci_master_dataa;             // NIOS_II_custom_instruction_master_translator:comb_ci_master_dataa -> NIOS_II_custom_instruction_master_comb_xconnect:ci_slave_dataa
	wire         nios_ii_custom_instruction_master_translator_comb_ci_master_writerc;           // NIOS_II_custom_instruction_master_translator:comb_ci_master_writerc -> NIOS_II_custom_instruction_master_comb_xconnect:ci_slave_writerc
	wire   [7:0] nios_ii_custom_instruction_master_translator_comb_ci_master_n;                 // NIOS_II_custom_instruction_master_translator:comb_ci_master_n -> NIOS_II_custom_instruction_master_comb_xconnect:ci_slave_n
	wire  [31:0] nios_ii_custom_instruction_master_comb_xconnect_ci_master0_result;             // NIOS_II_custom_instruction_master_comb_slave_translator0:ci_slave_result -> NIOS_II_custom_instruction_master_comb_xconnect:ci_master0_result
	wire         nios_ii_custom_instruction_master_comb_xconnect_ci_master0_readra;             // NIOS_II_custom_instruction_master_comb_xconnect:ci_master0_readra -> NIOS_II_custom_instruction_master_comb_slave_translator0:ci_slave_readra
	wire   [4:0] nios_ii_custom_instruction_master_comb_xconnect_ci_master0_a;                  // NIOS_II_custom_instruction_master_comb_xconnect:ci_master0_a -> NIOS_II_custom_instruction_master_comb_slave_translator0:ci_slave_a
	wire   [4:0] nios_ii_custom_instruction_master_comb_xconnect_ci_master0_b;                  // NIOS_II_custom_instruction_master_comb_xconnect:ci_master0_b -> NIOS_II_custom_instruction_master_comb_slave_translator0:ci_slave_b
	wire         nios_ii_custom_instruction_master_comb_xconnect_ci_master0_readrb;             // NIOS_II_custom_instruction_master_comb_xconnect:ci_master0_readrb -> NIOS_II_custom_instruction_master_comb_slave_translator0:ci_slave_readrb
	wire   [4:0] nios_ii_custom_instruction_master_comb_xconnect_ci_master0_c;                  // NIOS_II_custom_instruction_master_comb_xconnect:ci_master0_c -> NIOS_II_custom_instruction_master_comb_slave_translator0:ci_slave_c
	wire         nios_ii_custom_instruction_master_comb_xconnect_ci_master0_estatus;            // NIOS_II_custom_instruction_master_comb_xconnect:ci_master0_estatus -> NIOS_II_custom_instruction_master_comb_slave_translator0:ci_slave_estatus
	wire  [31:0] nios_ii_custom_instruction_master_comb_xconnect_ci_master0_ipending;           // NIOS_II_custom_instruction_master_comb_xconnect:ci_master0_ipending -> NIOS_II_custom_instruction_master_comb_slave_translator0:ci_slave_ipending
	wire  [31:0] nios_ii_custom_instruction_master_comb_xconnect_ci_master0_datab;              // NIOS_II_custom_instruction_master_comb_xconnect:ci_master0_datab -> NIOS_II_custom_instruction_master_comb_slave_translator0:ci_slave_datab
	wire  [31:0] nios_ii_custom_instruction_master_comb_xconnect_ci_master0_dataa;              // NIOS_II_custom_instruction_master_comb_xconnect:ci_master0_dataa -> NIOS_II_custom_instruction_master_comb_slave_translator0:ci_slave_dataa
	wire         nios_ii_custom_instruction_master_comb_xconnect_ci_master0_writerc;            // NIOS_II_custom_instruction_master_comb_xconnect:ci_master0_writerc -> NIOS_II_custom_instruction_master_comb_slave_translator0:ci_slave_writerc
	wire   [7:0] nios_ii_custom_instruction_master_comb_xconnect_ci_master0_n;                  // NIOS_II_custom_instruction_master_comb_xconnect:ci_master0_n -> NIOS_II_custom_instruction_master_comb_slave_translator0:ci_slave_n
	wire  [31:0] nios_ii_custom_instruction_master_comb_slave_translator0_ci_master_result;     // FPU:s1_result -> NIOS_II_custom_instruction_master_comb_slave_translator0:ci_master_result
	wire  [31:0] nios_ii_custom_instruction_master_comb_slave_translator0_ci_master_datab;      // NIOS_II_custom_instruction_master_comb_slave_translator0:ci_master_datab -> FPU:s1_datab
	wire  [31:0] nios_ii_custom_instruction_master_comb_slave_translator0_ci_master_dataa;      // NIOS_II_custom_instruction_master_comb_slave_translator0:ci_master_dataa -> FPU:s1_dataa
	wire   [3:0] nios_ii_custom_instruction_master_comb_slave_translator0_ci_master_n;          // NIOS_II_custom_instruction_master_comb_slave_translator0:ci_master_n -> FPU:s1_n
	wire         nios_ii_custom_instruction_master_translator_multi_ci_master_readra;           // NIOS_II_custom_instruction_master_translator:multi_ci_master_readra -> NIOS_II_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire   [4:0] nios_ii_custom_instruction_master_translator_multi_ci_master_a;                // NIOS_II_custom_instruction_master_translator:multi_ci_master_a -> NIOS_II_custom_instruction_master_multi_xconnect:ci_slave_a
	wire   [4:0] nios_ii_custom_instruction_master_translator_multi_ci_master_b;                // NIOS_II_custom_instruction_master_translator:multi_ci_master_b -> NIOS_II_custom_instruction_master_multi_xconnect:ci_slave_b
	wire         nios_ii_custom_instruction_master_translator_multi_ci_master_clk;              // NIOS_II_custom_instruction_master_translator:multi_ci_master_clk -> NIOS_II_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire         nios_ii_custom_instruction_master_translator_multi_ci_master_readrb;           // NIOS_II_custom_instruction_master_translator:multi_ci_master_readrb -> NIOS_II_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire   [4:0] nios_ii_custom_instruction_master_translator_multi_ci_master_c;                // NIOS_II_custom_instruction_master_translator:multi_ci_master_c -> NIOS_II_custom_instruction_master_multi_xconnect:ci_slave_c
	wire         nios_ii_custom_instruction_master_translator_multi_ci_master_start;            // NIOS_II_custom_instruction_master_translator:multi_ci_master_start -> NIOS_II_custom_instruction_master_multi_xconnect:ci_slave_start
	wire         nios_ii_custom_instruction_master_translator_multi_ci_master_reset_req;        // NIOS_II_custom_instruction_master_translator:multi_ci_master_reset_req -> NIOS_II_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	wire         nios_ii_custom_instruction_master_translator_multi_ci_master_done;             // NIOS_II_custom_instruction_master_multi_xconnect:ci_slave_done -> NIOS_II_custom_instruction_master_translator:multi_ci_master_done
	wire   [7:0] nios_ii_custom_instruction_master_translator_multi_ci_master_n;                // NIOS_II_custom_instruction_master_translator:multi_ci_master_n -> NIOS_II_custom_instruction_master_multi_xconnect:ci_slave_n
	wire  [31:0] nios_ii_custom_instruction_master_translator_multi_ci_master_result;           // NIOS_II_custom_instruction_master_multi_xconnect:ci_slave_result -> NIOS_II_custom_instruction_master_translator:multi_ci_master_result
	wire         nios_ii_custom_instruction_master_translator_multi_ci_master_clk_en;           // NIOS_II_custom_instruction_master_translator:multi_ci_master_clken -> NIOS_II_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire  [31:0] nios_ii_custom_instruction_master_translator_multi_ci_master_datab;            // NIOS_II_custom_instruction_master_translator:multi_ci_master_datab -> NIOS_II_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire  [31:0] nios_ii_custom_instruction_master_translator_multi_ci_master_dataa;            // NIOS_II_custom_instruction_master_translator:multi_ci_master_dataa -> NIOS_II_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire         nios_ii_custom_instruction_master_translator_multi_ci_master_reset;            // NIOS_II_custom_instruction_master_translator:multi_ci_master_reset -> NIOS_II_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire         nios_ii_custom_instruction_master_translator_multi_ci_master_writerc;          // NIOS_II_custom_instruction_master_translator:multi_ci_master_writerc -> NIOS_II_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire         nios_ii_custom_instruction_master_multi_xconnect_ci_master0_readra;            // NIOS_II_custom_instruction_master_multi_xconnect:ci_master0_readra -> NIOS_II_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire   [4:0] nios_ii_custom_instruction_master_multi_xconnect_ci_master0_a;                 // NIOS_II_custom_instruction_master_multi_xconnect:ci_master0_a -> NIOS_II_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire   [4:0] nios_ii_custom_instruction_master_multi_xconnect_ci_master0_b;                 // NIOS_II_custom_instruction_master_multi_xconnect:ci_master0_b -> NIOS_II_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire         nios_ii_custom_instruction_master_multi_xconnect_ci_master0_readrb;            // NIOS_II_custom_instruction_master_multi_xconnect:ci_master0_readrb -> NIOS_II_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire   [4:0] nios_ii_custom_instruction_master_multi_xconnect_ci_master0_c;                 // NIOS_II_custom_instruction_master_multi_xconnect:ci_master0_c -> NIOS_II_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire         nios_ii_custom_instruction_master_multi_xconnect_ci_master0_clk;               // NIOS_II_custom_instruction_master_multi_xconnect:ci_master0_clk -> NIOS_II_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire  [31:0] nios_ii_custom_instruction_master_multi_xconnect_ci_master0_ipending;          // NIOS_II_custom_instruction_master_multi_xconnect:ci_master0_ipending -> NIOS_II_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire         nios_ii_custom_instruction_master_multi_xconnect_ci_master0_start;             // NIOS_II_custom_instruction_master_multi_xconnect:ci_master0_start -> NIOS_II_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire         nios_ii_custom_instruction_master_multi_xconnect_ci_master0_reset_req;         // NIOS_II_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> NIOS_II_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	wire         nios_ii_custom_instruction_master_multi_xconnect_ci_master0_done;              // NIOS_II_custom_instruction_master_multi_slave_translator0:ci_slave_done -> NIOS_II_custom_instruction_master_multi_xconnect:ci_master0_done
	wire   [7:0] nios_ii_custom_instruction_master_multi_xconnect_ci_master0_n;                 // NIOS_II_custom_instruction_master_multi_xconnect:ci_master0_n -> NIOS_II_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire  [31:0] nios_ii_custom_instruction_master_multi_xconnect_ci_master0_result;            // NIOS_II_custom_instruction_master_multi_slave_translator0:ci_slave_result -> NIOS_II_custom_instruction_master_multi_xconnect:ci_master0_result
	wire         nios_ii_custom_instruction_master_multi_xconnect_ci_master0_estatus;           // NIOS_II_custom_instruction_master_multi_xconnect:ci_master0_estatus -> NIOS_II_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire         nios_ii_custom_instruction_master_multi_xconnect_ci_master0_clk_en;            // NIOS_II_custom_instruction_master_multi_xconnect:ci_master0_clken -> NIOS_II_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire  [31:0] nios_ii_custom_instruction_master_multi_xconnect_ci_master0_datab;             // NIOS_II_custom_instruction_master_multi_xconnect:ci_master0_datab -> NIOS_II_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire  [31:0] nios_ii_custom_instruction_master_multi_xconnect_ci_master0_dataa;             // NIOS_II_custom_instruction_master_multi_xconnect:ci_master0_dataa -> NIOS_II_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire         nios_ii_custom_instruction_master_multi_xconnect_ci_master0_reset;             // NIOS_II_custom_instruction_master_multi_xconnect:ci_master0_reset -> NIOS_II_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire         nios_ii_custom_instruction_master_multi_xconnect_ci_master0_writerc;           // NIOS_II_custom_instruction_master_multi_xconnect:ci_master0_writerc -> NIOS_II_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire  [31:0] nios_ii_custom_instruction_master_multi_slave_translator0_ci_master_result;    // FPU:s2_result -> NIOS_II_custom_instruction_master_multi_slave_translator0:ci_master_result
	wire         nios_ii_custom_instruction_master_multi_slave_translator0_ci_master_clk;       // NIOS_II_custom_instruction_master_multi_slave_translator0:ci_master_clk -> FPU:s2_clk
	wire         nios_ii_custom_instruction_master_multi_slave_translator0_ci_master_clk_en;    // NIOS_II_custom_instruction_master_multi_slave_translator0:ci_master_clken -> FPU:s2_clk_en
	wire  [31:0] nios_ii_custom_instruction_master_multi_slave_translator0_ci_master_datab;     // NIOS_II_custom_instruction_master_multi_slave_translator0:ci_master_datab -> FPU:s2_datab
	wire  [31:0] nios_ii_custom_instruction_master_multi_slave_translator0_ci_master_dataa;     // NIOS_II_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> FPU:s2_dataa
	wire         nios_ii_custom_instruction_master_multi_slave_translator0_ci_master_start;     // NIOS_II_custom_instruction_master_multi_slave_translator0:ci_master_start -> FPU:s2_start
	wire         nios_ii_custom_instruction_master_multi_slave_translator0_ci_master_reset;     // NIOS_II_custom_instruction_master_multi_slave_translator0:ci_master_reset -> FPU:s2_reset
	wire         nios_ii_custom_instruction_master_multi_slave_translator0_ci_master_reset_req; // NIOS_II_custom_instruction_master_multi_slave_translator0:ci_master_reset_req -> FPU:s2_reset_req
	wire         nios_ii_custom_instruction_master_multi_slave_translator0_ci_master_done;      // FPU:s2_done -> NIOS_II_custom_instruction_master_multi_slave_translator0:ci_master_done
	wire   [2:0] nios_ii_custom_instruction_master_multi_slave_translator0_ci_master_n;         // NIOS_II_custom_instruction_master_multi_slave_translator0:ci_master_n -> FPU:s2_n
	wire  [31:0] nios_ii_data_master_readdata;                                                  // mm_interconnect_0:NIOS_II_data_master_readdata -> NIOS_II:d_readdata
	wire         nios_ii_data_master_waitrequest;                                               // mm_interconnect_0:NIOS_II_data_master_waitrequest -> NIOS_II:d_waitrequest
	wire         nios_ii_data_master_debugaccess;                                               // NIOS_II:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NIOS_II_data_master_debugaccess
	wire  [19:0] nios_ii_data_master_address;                                                   // NIOS_II:d_address -> mm_interconnect_0:NIOS_II_data_master_address
	wire   [3:0] nios_ii_data_master_byteenable;                                                // NIOS_II:d_byteenable -> mm_interconnect_0:NIOS_II_data_master_byteenable
	wire         nios_ii_data_master_read;                                                      // NIOS_II:d_read -> mm_interconnect_0:NIOS_II_data_master_read
	wire         nios_ii_data_master_write;                                                     // NIOS_II:d_write -> mm_interconnect_0:NIOS_II_data_master_write
	wire  [31:0] nios_ii_data_master_writedata;                                                 // NIOS_II:d_writedata -> mm_interconnect_0:NIOS_II_data_master_writedata
	wire  [31:0] nios_ii_instruction_master_readdata;                                           // mm_interconnect_0:NIOS_II_instruction_master_readdata -> NIOS_II:i_readdata
	wire         nios_ii_instruction_master_waitrequest;                                        // mm_interconnect_0:NIOS_II_instruction_master_waitrequest -> NIOS_II:i_waitrequest
	wire  [19:0] nios_ii_instruction_master_address;                                            // NIOS_II:i_address -> mm_interconnect_0:NIOS_II_instruction_master_address
	wire         nios_ii_instruction_master_read;                                               // NIOS_II:i_read -> mm_interconnect_0:NIOS_II_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;                      // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_chipselect -> JTAG_UART:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;                        // JTAG_UART:av_readdata -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;                     // JTAG_UART:av_waitrequest -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;                         // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_address -> JTAG_UART:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                            // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_read -> JTAG_UART:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                           // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_write -> JTAG_UART:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;                       // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_writedata -> JTAG_UART:av_writedata
	wire  [31:0] mm_interconnect_0_performance_counter_control_slave_readdata;                  // PERFORMANCE_COUNTER:readdata -> mm_interconnect_0:PERFORMANCE_COUNTER_control_slave_readdata
	wire   [3:0] mm_interconnect_0_performance_counter_control_slave_address;                   // mm_interconnect_0:PERFORMANCE_COUNTER_control_slave_address -> PERFORMANCE_COUNTER:address
	wire         mm_interconnect_0_performance_counter_control_slave_begintransfer;             // mm_interconnect_0:PERFORMANCE_COUNTER_control_slave_begintransfer -> PERFORMANCE_COUNTER:begintransfer
	wire         mm_interconnect_0_performance_counter_control_slave_write;                     // mm_interconnect_0:PERFORMANCE_COUNTER_control_slave_write -> PERFORMANCE_COUNTER:write
	wire  [31:0] mm_interconnect_0_performance_counter_control_slave_writedata;                 // mm_interconnect_0:PERFORMANCE_COUNTER_control_slave_writedata -> PERFORMANCE_COUNTER:writedata
	wire  [31:0] mm_interconnect_0_nios_ii_debug_mem_slave_readdata;                            // NIOS_II:debug_mem_slave_readdata -> mm_interconnect_0:NIOS_II_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios_ii_debug_mem_slave_waitrequest;                         // NIOS_II:debug_mem_slave_waitrequest -> mm_interconnect_0:NIOS_II_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios_ii_debug_mem_slave_debugaccess;                         // mm_interconnect_0:NIOS_II_debug_mem_slave_debugaccess -> NIOS_II:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios_ii_debug_mem_slave_address;                             // mm_interconnect_0:NIOS_II_debug_mem_slave_address -> NIOS_II:debug_mem_slave_address
	wire         mm_interconnect_0_nios_ii_debug_mem_slave_read;                                // mm_interconnect_0:NIOS_II_debug_mem_slave_read -> NIOS_II:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios_ii_debug_mem_slave_byteenable;                          // mm_interconnect_0:NIOS_II_debug_mem_slave_byteenable -> NIOS_II:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios_ii_debug_mem_slave_write;                               // mm_interconnect_0:NIOS_II_debug_mem_slave_write -> NIOS_II:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios_ii_debug_mem_slave_writedata;                           // mm_interconnect_0:NIOS_II_debug_mem_slave_writedata -> NIOS_II:debug_mem_slave_writedata
	wire         mm_interconnect_0_ram_s1_chipselect;                                           // mm_interconnect_0:RAM_s1_chipselect -> RAM:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                                             // RAM:readdata -> mm_interconnect_0:RAM_s1_readdata
	wire  [15:0] mm_interconnect_0_ram_s1_address;                                              // mm_interconnect_0:RAM_s1_address -> RAM:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;                                           // mm_interconnect_0:RAM_s1_byteenable -> RAM:byteenable
	wire         mm_interconnect_0_ram_s1_write;                                                // mm_interconnect_0:RAM_s1_write -> RAM:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                                            // mm_interconnect_0:RAM_s1_writedata -> RAM:writedata
	wire         mm_interconnect_0_ram_s1_clken;                                                // mm_interconnect_0:RAM_s1_clken -> RAM:clken
	wire         irq_mapper_receiver0_irq;                                                      // JTAG_UART:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios_ii_irq_irq;                                                               // irq_mapper:sender_irq -> NIOS_II:irq
	wire         rst_controller_reset_out_reset;                                                // rst_controller:reset_out -> [JTAG_UART:rst_n, NIOS_II:reset_n, PERFORMANCE_COUNTER:reset_n, RAM:reset, irq_mapper:reset, mm_interconnect_0:NIOS_II_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                                            // rst_controller:reset_req -> [NIOS_II:reset_req, RAM:reset_req, rst_translator:reset_req_in]
	wire         nios_ii_debug_reset_request_reset;                                             // NIOS_II:debug_reset_request -> rst_controller:reset_in1

	Nios2_accelerator_FPU #(
		.arithmetic_present (1),
		.root_present       (0),
		.conversion_present (1),
		.comparison_present (0)
	) fpu (
		.s1_dataa     (nios_ii_custom_instruction_master_comb_slave_translator0_ci_master_dataa),      // s1.dataa
		.s1_datab     (nios_ii_custom_instruction_master_comb_slave_translator0_ci_master_datab),      //   .datab
		.s1_n         (nios_ii_custom_instruction_master_comb_slave_translator0_ci_master_n),          //   .n
		.s1_result    (nios_ii_custom_instruction_master_comb_slave_translator0_ci_master_result),     //   .result
		.s2_clk       (nios_ii_custom_instruction_master_multi_slave_translator0_ci_master_clk),       // s2.clk
		.s2_clk_en    (nios_ii_custom_instruction_master_multi_slave_translator0_ci_master_clk_en),    //   .clk_en
		.s2_dataa     (nios_ii_custom_instruction_master_multi_slave_translator0_ci_master_dataa),     //   .dataa
		.s2_datab     (nios_ii_custom_instruction_master_multi_slave_translator0_ci_master_datab),     //   .datab
		.s2_n         (nios_ii_custom_instruction_master_multi_slave_translator0_ci_master_n),         //   .n
		.s2_reset     (nios_ii_custom_instruction_master_multi_slave_translator0_ci_master_reset),     //   .reset
		.s2_reset_req (nios_ii_custom_instruction_master_multi_slave_translator0_ci_master_reset_req), //   .reset_req
		.s2_start     (nios_ii_custom_instruction_master_multi_slave_translator0_ci_master_start),     //   .start
		.s2_done      (nios_ii_custom_instruction_master_multi_slave_translator0_ci_master_done),      //   .done
		.s2_result    (nios_ii_custom_instruction_master_multi_slave_translator0_ci_master_result)     //   .result
	);

	Nios2_accelerator_JTAG_UART jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	Nios2_accelerator_NIOS_II nios_ii (
		.clk                                 (clk_clk),                                               //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                       //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                    //                          .reset_req
		.d_address                           (nios_ii_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios_ii_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios_ii_data_master_read),                              //                          .read
		.d_readdata                          (nios_ii_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios_ii_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios_ii_data_master_write),                             //                          .write
		.d_writedata                         (nios_ii_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios_ii_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios_ii_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios_ii_instruction_master_read),                       //                          .read
		.i_readdata                          (nios_ii_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios_ii_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios_ii_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios_ii_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios_ii_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios_ii_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios_ii_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios_ii_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios_ii_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios_ii_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios_ii_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios_ii_debug_mem_slave_writedata),   //                          .writedata
		.E_ci_multi_done                     (nios_ii_custom_instruction_master_done),                // custom_instruction_master.done
		.E_ci_multi_clk_en                   (nios_ii_custom_instruction_master_clk_en),              //                          .clk_en
		.E_ci_multi_start                    (nios_ii_custom_instruction_master_start),               //                          .start
		.E_ci_result                         (nios_ii_custom_instruction_master_result),              //                          .result
		.D_ci_a                              (nios_ii_custom_instruction_master_a),                   //                          .a
		.D_ci_b                              (nios_ii_custom_instruction_master_b),                   //                          .b
		.D_ci_c                              (nios_ii_custom_instruction_master_c),                   //                          .c
		.D_ci_n                              (nios_ii_custom_instruction_master_n),                   //                          .n
		.D_ci_readra                         (nios_ii_custom_instruction_master_readra),              //                          .readra
		.D_ci_readrb                         (nios_ii_custom_instruction_master_readrb),              //                          .readrb
		.D_ci_writerc                        (nios_ii_custom_instruction_master_writerc),             //                          .writerc
		.E_ci_dataa                          (nios_ii_custom_instruction_master_dataa),               //                          .dataa
		.E_ci_datab                          (nios_ii_custom_instruction_master_datab),               //                          .datab
		.E_ci_multi_clock                    (nios_ii_custom_instruction_master_clk),                 //                          .clk
		.E_ci_multi_reset                    (nios_ii_custom_instruction_master_reset),               //                          .reset
		.E_ci_multi_reset_req                (nios_ii_custom_instruction_master_reset_req),           //                          .reset_req
		.W_ci_estatus                        (nios_ii_custom_instruction_master_estatus),             //                          .estatus
		.W_ci_ipending                       (nios_ii_custom_instruction_master_ipending)             //                          .ipending
	);

	Nios2_accelerator_PERFORMANCE_COUNTER performance_counter (
		.clk           (clk_clk),                                                           //           clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                                   //         reset.reset_n
		.address       (mm_interconnect_0_performance_counter_control_slave_address),       // control_slave.address
		.begintransfer (mm_interconnect_0_performance_counter_control_slave_begintransfer), //              .begintransfer
		.readdata      (mm_interconnect_0_performance_counter_control_slave_readdata),      //              .readdata
		.write         (mm_interconnect_0_performance_counter_control_slave_write),         //              .write
		.writedata     (mm_interconnect_0_performance_counter_control_slave_writedata)      //              .writedata
	);

	Nios2_accelerator_RAM ram (
		.clk        (clk_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze     (1'b0)                                 // (terminated)
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (1)
	) nios_ii_custom_instruction_master_translator (
		.ci_slave_dataa            (nios_ii_custom_instruction_master_dataa),                                //        ci_slave.dataa
		.ci_slave_datab            (nios_ii_custom_instruction_master_datab),                                //                .datab
		.ci_slave_result           (nios_ii_custom_instruction_master_result),                               //                .result
		.ci_slave_n                (nios_ii_custom_instruction_master_n),                                    //                .n
		.ci_slave_readra           (nios_ii_custom_instruction_master_readra),                               //                .readra
		.ci_slave_readrb           (nios_ii_custom_instruction_master_readrb),                               //                .readrb
		.ci_slave_writerc          (nios_ii_custom_instruction_master_writerc),                              //                .writerc
		.ci_slave_a                (nios_ii_custom_instruction_master_a),                                    //                .a
		.ci_slave_b                (nios_ii_custom_instruction_master_b),                                    //                .b
		.ci_slave_c                (nios_ii_custom_instruction_master_c),                                    //                .c
		.ci_slave_ipending         (nios_ii_custom_instruction_master_ipending),                             //                .ipending
		.ci_slave_estatus          (nios_ii_custom_instruction_master_estatus),                              //                .estatus
		.ci_slave_multi_clk        (nios_ii_custom_instruction_master_clk),                                  //                .clk
		.ci_slave_multi_reset      (nios_ii_custom_instruction_master_reset),                                //                .reset
		.ci_slave_multi_clken      (nios_ii_custom_instruction_master_clk_en),                               //                .clk_en
		.ci_slave_multi_reset_req  (nios_ii_custom_instruction_master_reset_req),                            //                .reset_req
		.ci_slave_multi_start      (nios_ii_custom_instruction_master_start),                                //                .start
		.ci_slave_multi_done       (nios_ii_custom_instruction_master_done),                                 //                .done
		.comb_ci_master_dataa      (nios_ii_custom_instruction_master_translator_comb_ci_master_dataa),      //  comb_ci_master.dataa
		.comb_ci_master_datab      (nios_ii_custom_instruction_master_translator_comb_ci_master_datab),      //                .datab
		.comb_ci_master_result     (nios_ii_custom_instruction_master_translator_comb_ci_master_result),     //                .result
		.comb_ci_master_n          (nios_ii_custom_instruction_master_translator_comb_ci_master_n),          //                .n
		.comb_ci_master_readra     (nios_ii_custom_instruction_master_translator_comb_ci_master_readra),     //                .readra
		.comb_ci_master_readrb     (nios_ii_custom_instruction_master_translator_comb_ci_master_readrb),     //                .readrb
		.comb_ci_master_writerc    (nios_ii_custom_instruction_master_translator_comb_ci_master_writerc),    //                .writerc
		.comb_ci_master_a          (nios_ii_custom_instruction_master_translator_comb_ci_master_a),          //                .a
		.comb_ci_master_b          (nios_ii_custom_instruction_master_translator_comb_ci_master_b),          //                .b
		.comb_ci_master_c          (nios_ii_custom_instruction_master_translator_comb_ci_master_c),          //                .c
		.comb_ci_master_ipending   (nios_ii_custom_instruction_master_translator_comb_ci_master_ipending),   //                .ipending
		.comb_ci_master_estatus    (nios_ii_custom_instruction_master_translator_comb_ci_master_estatus),    //                .estatus
		.multi_ci_master_clk       (nios_ii_custom_instruction_master_translator_multi_ci_master_clk),       // multi_ci_master.clk
		.multi_ci_master_reset     (nios_ii_custom_instruction_master_translator_multi_ci_master_reset),     //                .reset
		.multi_ci_master_clken     (nios_ii_custom_instruction_master_translator_multi_ci_master_clk_en),    //                .clk_en
		.multi_ci_master_reset_req (nios_ii_custom_instruction_master_translator_multi_ci_master_reset_req), //                .reset_req
		.multi_ci_master_start     (nios_ii_custom_instruction_master_translator_multi_ci_master_start),     //                .start
		.multi_ci_master_done      (nios_ii_custom_instruction_master_translator_multi_ci_master_done),      //                .done
		.multi_ci_master_dataa     (nios_ii_custom_instruction_master_translator_multi_ci_master_dataa),     //                .dataa
		.multi_ci_master_datab     (nios_ii_custom_instruction_master_translator_multi_ci_master_datab),     //                .datab
		.multi_ci_master_result    (nios_ii_custom_instruction_master_translator_multi_ci_master_result),    //                .result
		.multi_ci_master_n         (nios_ii_custom_instruction_master_translator_multi_ci_master_n),         //                .n
		.multi_ci_master_readra    (nios_ii_custom_instruction_master_translator_multi_ci_master_readra),    //                .readra
		.multi_ci_master_readrb    (nios_ii_custom_instruction_master_translator_multi_ci_master_readrb),    //                .readrb
		.multi_ci_master_writerc   (nios_ii_custom_instruction_master_translator_multi_ci_master_writerc),   //                .writerc
		.multi_ci_master_a         (nios_ii_custom_instruction_master_translator_multi_ci_master_a),         //                .a
		.multi_ci_master_b         (nios_ii_custom_instruction_master_translator_multi_ci_master_b),         //                .b
		.multi_ci_master_c         (nios_ii_custom_instruction_master_translator_multi_ci_master_c),         //                .c
		.ci_slave_multi_dataa      (32'b00000000000000000000000000000000),                                   //     (terminated)
		.ci_slave_multi_datab      (32'b00000000000000000000000000000000),                                   //     (terminated)
		.ci_slave_multi_result     (),                                                                       //     (terminated)
		.ci_slave_multi_n          (8'b00000000),                                                            //     (terminated)
		.ci_slave_multi_readra     (1'b0),                                                                   //     (terminated)
		.ci_slave_multi_readrb     (1'b0),                                                                   //     (terminated)
		.ci_slave_multi_writerc    (1'b0),                                                                   //     (terminated)
		.ci_slave_multi_a          (5'b00000),                                                               //     (terminated)
		.ci_slave_multi_b          (5'b00000),                                                               //     (terminated)
		.ci_slave_multi_c          (5'b00000)                                                                //     (terminated)
	);

	Nios2_accelerator_NIOS_II_custom_instruction_master_comb_xconnect nios_ii_custom_instruction_master_comb_xconnect (
		.ci_slave_dataa      (nios_ii_custom_instruction_master_translator_comb_ci_master_dataa),    //   ci_slave.dataa
		.ci_slave_datab      (nios_ii_custom_instruction_master_translator_comb_ci_master_datab),    //           .datab
		.ci_slave_result     (nios_ii_custom_instruction_master_translator_comb_ci_master_result),   //           .result
		.ci_slave_n          (nios_ii_custom_instruction_master_translator_comb_ci_master_n),        //           .n
		.ci_slave_readra     (nios_ii_custom_instruction_master_translator_comb_ci_master_readra),   //           .readra
		.ci_slave_readrb     (nios_ii_custom_instruction_master_translator_comb_ci_master_readrb),   //           .readrb
		.ci_slave_writerc    (nios_ii_custom_instruction_master_translator_comb_ci_master_writerc),  //           .writerc
		.ci_slave_a          (nios_ii_custom_instruction_master_translator_comb_ci_master_a),        //           .a
		.ci_slave_b          (nios_ii_custom_instruction_master_translator_comb_ci_master_b),        //           .b
		.ci_slave_c          (nios_ii_custom_instruction_master_translator_comb_ci_master_c),        //           .c
		.ci_slave_ipending   (nios_ii_custom_instruction_master_translator_comb_ci_master_ipending), //           .ipending
		.ci_slave_estatus    (nios_ii_custom_instruction_master_translator_comb_ci_master_estatus),  //           .estatus
		.ci_master0_dataa    (nios_ii_custom_instruction_master_comb_xconnect_ci_master0_dataa),     // ci_master0.dataa
		.ci_master0_datab    (nios_ii_custom_instruction_master_comb_xconnect_ci_master0_datab),     //           .datab
		.ci_master0_result   (nios_ii_custom_instruction_master_comb_xconnect_ci_master0_result),    //           .result
		.ci_master0_n        (nios_ii_custom_instruction_master_comb_xconnect_ci_master0_n),         //           .n
		.ci_master0_readra   (nios_ii_custom_instruction_master_comb_xconnect_ci_master0_readra),    //           .readra
		.ci_master0_readrb   (nios_ii_custom_instruction_master_comb_xconnect_ci_master0_readrb),    //           .readrb
		.ci_master0_writerc  (nios_ii_custom_instruction_master_comb_xconnect_ci_master0_writerc),   //           .writerc
		.ci_master0_a        (nios_ii_custom_instruction_master_comb_xconnect_ci_master0_a),         //           .a
		.ci_master0_b        (nios_ii_custom_instruction_master_comb_xconnect_ci_master0_b),         //           .b
		.ci_master0_c        (nios_ii_custom_instruction_master_comb_xconnect_ci_master0_c),         //           .c
		.ci_master0_ipending (nios_ii_custom_instruction_master_comb_xconnect_ci_master0_ipending),  //           .ipending
		.ci_master0_estatus  (nios_ii_custom_instruction_master_comb_xconnect_ci_master0_estatus)    //           .estatus
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (4),
		.USE_DONE         (0),
		.NUM_FIXED_CYCLES (0)
	) nios_ii_custom_instruction_master_comb_slave_translator0 (
		.ci_slave_dataa      (nios_ii_custom_instruction_master_comb_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios_ii_custom_instruction_master_comb_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (nios_ii_custom_instruction_master_comb_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (nios_ii_custom_instruction_master_comb_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (nios_ii_custom_instruction_master_comb_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (nios_ii_custom_instruction_master_comb_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (nios_ii_custom_instruction_master_comb_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (nios_ii_custom_instruction_master_comb_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (nios_ii_custom_instruction_master_comb_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (nios_ii_custom_instruction_master_comb_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (nios_ii_custom_instruction_master_comb_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (nios_ii_custom_instruction_master_comb_xconnect_ci_master0_estatus),        //          .estatus
		.ci_master_dataa     (nios_ii_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios_ii_custom_instruction_master_comb_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (nios_ii_custom_instruction_master_comb_slave_translator0_ci_master_result), //          .result
		.ci_master_n         (nios_ii_custom_instruction_master_comb_slave_translator0_ci_master_n),      //          .n
		.ci_master_readra    (),                                                                          // (terminated)
		.ci_master_readrb    (),                                                                          // (terminated)
		.ci_master_writerc   (),                                                                          // (terminated)
		.ci_master_a         (),                                                                          // (terminated)
		.ci_master_b         (),                                                                          // (terminated)
		.ci_master_c         (),                                                                          // (terminated)
		.ci_master_ipending  (),                                                                          // (terminated)
		.ci_master_estatus   (),                                                                          // (terminated)
		.ci_master_clk       (),                                                                          // (terminated)
		.ci_master_clken     (),                                                                          // (terminated)
		.ci_master_reset_req (),                                                                          // (terminated)
		.ci_master_reset     (),                                                                          // (terminated)
		.ci_master_start     (),                                                                          // (terminated)
		.ci_master_done      (1'b0),                                                                      // (terminated)
		.ci_slave_clk        (1'b0),                                                                      // (terminated)
		.ci_slave_clken      (1'b0),                                                                      // (terminated)
		.ci_slave_reset_req  (1'b0),                                                                      // (terminated)
		.ci_slave_reset      (1'b0),                                                                      // (terminated)
		.ci_slave_start      (1'b0),                                                                      // (terminated)
		.ci_slave_done       ()                                                                           // (terminated)
	);

	Nios2_accelerator_NIOS_II_custom_instruction_master_multi_xconnect nios_ii_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa       (nios_ii_custom_instruction_master_translator_multi_ci_master_dataa),     //   ci_slave.dataa
		.ci_slave_datab       (nios_ii_custom_instruction_master_translator_multi_ci_master_datab),     //           .datab
		.ci_slave_result      (nios_ii_custom_instruction_master_translator_multi_ci_master_result),    //           .result
		.ci_slave_n           (nios_ii_custom_instruction_master_translator_multi_ci_master_n),         //           .n
		.ci_slave_readra      (nios_ii_custom_instruction_master_translator_multi_ci_master_readra),    //           .readra
		.ci_slave_readrb      (nios_ii_custom_instruction_master_translator_multi_ci_master_readrb),    //           .readrb
		.ci_slave_writerc     (nios_ii_custom_instruction_master_translator_multi_ci_master_writerc),   //           .writerc
		.ci_slave_a           (nios_ii_custom_instruction_master_translator_multi_ci_master_a),         //           .a
		.ci_slave_b           (nios_ii_custom_instruction_master_translator_multi_ci_master_b),         //           .b
		.ci_slave_c           (nios_ii_custom_instruction_master_translator_multi_ci_master_c),         //           .c
		.ci_slave_ipending    (),                                                                       //           .ipending
		.ci_slave_estatus     (),                                                                       //           .estatus
		.ci_slave_clk         (nios_ii_custom_instruction_master_translator_multi_ci_master_clk),       //           .clk
		.ci_slave_reset       (nios_ii_custom_instruction_master_translator_multi_ci_master_reset),     //           .reset
		.ci_slave_clken       (nios_ii_custom_instruction_master_translator_multi_ci_master_clk_en),    //           .clk_en
		.ci_slave_reset_req   (nios_ii_custom_instruction_master_translator_multi_ci_master_reset_req), //           .reset_req
		.ci_slave_start       (nios_ii_custom_instruction_master_translator_multi_ci_master_start),     //           .start
		.ci_slave_done        (nios_ii_custom_instruction_master_translator_multi_ci_master_done),      //           .done
		.ci_master0_dataa     (nios_ii_custom_instruction_master_multi_xconnect_ci_master0_dataa),      // ci_master0.dataa
		.ci_master0_datab     (nios_ii_custom_instruction_master_multi_xconnect_ci_master0_datab),      //           .datab
		.ci_master0_result    (nios_ii_custom_instruction_master_multi_xconnect_ci_master0_result),     //           .result
		.ci_master0_n         (nios_ii_custom_instruction_master_multi_xconnect_ci_master0_n),          //           .n
		.ci_master0_readra    (nios_ii_custom_instruction_master_multi_xconnect_ci_master0_readra),     //           .readra
		.ci_master0_readrb    (nios_ii_custom_instruction_master_multi_xconnect_ci_master0_readrb),     //           .readrb
		.ci_master0_writerc   (nios_ii_custom_instruction_master_multi_xconnect_ci_master0_writerc),    //           .writerc
		.ci_master0_a         (nios_ii_custom_instruction_master_multi_xconnect_ci_master0_a),          //           .a
		.ci_master0_b         (nios_ii_custom_instruction_master_multi_xconnect_ci_master0_b),          //           .b
		.ci_master0_c         (nios_ii_custom_instruction_master_multi_xconnect_ci_master0_c),          //           .c
		.ci_master0_ipending  (nios_ii_custom_instruction_master_multi_xconnect_ci_master0_ipending),   //           .ipending
		.ci_master0_estatus   (nios_ii_custom_instruction_master_multi_xconnect_ci_master0_estatus),    //           .estatus
		.ci_master0_clk       (nios_ii_custom_instruction_master_multi_xconnect_ci_master0_clk),        //           .clk
		.ci_master0_reset     (nios_ii_custom_instruction_master_multi_xconnect_ci_master0_reset),      //           .reset
		.ci_master0_clken     (nios_ii_custom_instruction_master_multi_xconnect_ci_master0_clk_en),     //           .clk_en
		.ci_master0_reset_req (nios_ii_custom_instruction_master_multi_xconnect_ci_master0_reset_req),  //           .reset_req
		.ci_master0_start     (nios_ii_custom_instruction_master_multi_xconnect_ci_master0_start),      //           .start
		.ci_master0_done      (nios_ii_custom_instruction_master_multi_xconnect_ci_master0_done)        //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (3),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (1)
	) nios_ii_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa      (nios_ii_custom_instruction_master_multi_xconnect_ci_master0_dataa),             //  ci_slave.dataa
		.ci_slave_datab      (nios_ii_custom_instruction_master_multi_xconnect_ci_master0_datab),             //          .datab
		.ci_slave_result     (nios_ii_custom_instruction_master_multi_xconnect_ci_master0_result),            //          .result
		.ci_slave_n          (nios_ii_custom_instruction_master_multi_xconnect_ci_master0_n),                 //          .n
		.ci_slave_readra     (nios_ii_custom_instruction_master_multi_xconnect_ci_master0_readra),            //          .readra
		.ci_slave_readrb     (nios_ii_custom_instruction_master_multi_xconnect_ci_master0_readrb),            //          .readrb
		.ci_slave_writerc    (nios_ii_custom_instruction_master_multi_xconnect_ci_master0_writerc),           //          .writerc
		.ci_slave_a          (nios_ii_custom_instruction_master_multi_xconnect_ci_master0_a),                 //          .a
		.ci_slave_b          (nios_ii_custom_instruction_master_multi_xconnect_ci_master0_b),                 //          .b
		.ci_slave_c          (nios_ii_custom_instruction_master_multi_xconnect_ci_master0_c),                 //          .c
		.ci_slave_ipending   (nios_ii_custom_instruction_master_multi_xconnect_ci_master0_ipending),          //          .ipending
		.ci_slave_estatus    (nios_ii_custom_instruction_master_multi_xconnect_ci_master0_estatus),           //          .estatus
		.ci_slave_clk        (nios_ii_custom_instruction_master_multi_xconnect_ci_master0_clk),               //          .clk
		.ci_slave_clken      (nios_ii_custom_instruction_master_multi_xconnect_ci_master0_clk_en),            //          .clk_en
		.ci_slave_reset_req  (nios_ii_custom_instruction_master_multi_xconnect_ci_master0_reset_req),         //          .reset_req
		.ci_slave_reset      (nios_ii_custom_instruction_master_multi_xconnect_ci_master0_reset),             //          .reset
		.ci_slave_start      (nios_ii_custom_instruction_master_multi_xconnect_ci_master0_start),             //          .start
		.ci_slave_done       (nios_ii_custom_instruction_master_multi_xconnect_ci_master0_done),              //          .done
		.ci_master_dataa     (nios_ii_custom_instruction_master_multi_slave_translator0_ci_master_dataa),     // ci_master.dataa
		.ci_master_datab     (nios_ii_custom_instruction_master_multi_slave_translator0_ci_master_datab),     //          .datab
		.ci_master_result    (nios_ii_custom_instruction_master_multi_slave_translator0_ci_master_result),    //          .result
		.ci_master_n         (nios_ii_custom_instruction_master_multi_slave_translator0_ci_master_n),         //          .n
		.ci_master_clk       (nios_ii_custom_instruction_master_multi_slave_translator0_ci_master_clk),       //          .clk
		.ci_master_clken     (nios_ii_custom_instruction_master_multi_slave_translator0_ci_master_clk_en),    //          .clk_en
		.ci_master_reset_req (nios_ii_custom_instruction_master_multi_slave_translator0_ci_master_reset_req), //          .reset_req
		.ci_master_reset     (nios_ii_custom_instruction_master_multi_slave_translator0_ci_master_reset),     //          .reset
		.ci_master_start     (nios_ii_custom_instruction_master_multi_slave_translator0_ci_master_start),     //          .start
		.ci_master_done      (nios_ii_custom_instruction_master_multi_slave_translator0_ci_master_done),      //          .done
		.ci_master_readra    (),                                                                              // (terminated)
		.ci_master_readrb    (),                                                                              // (terminated)
		.ci_master_writerc   (),                                                                              // (terminated)
		.ci_master_a         (),                                                                              // (terminated)
		.ci_master_b         (),                                                                              // (terminated)
		.ci_master_c         (),                                                                              // (terminated)
		.ci_master_ipending  (),                                                                              // (terminated)
		.ci_master_estatus   ()                                                                               // (terminated)
	);

	Nios2_accelerator_mm_interconnect_0 mm_interconnect_0 (
		.CLK_clk_clk                                     (clk_clk),                                                           //                             CLK_clk.clk
		.NIOS_II_reset_reset_bridge_in_reset_reset       (rst_controller_reset_out_reset),                                    // NIOS_II_reset_reset_bridge_in_reset.reset
		.NIOS_II_data_master_address                     (nios_ii_data_master_address),                                       //                 NIOS_II_data_master.address
		.NIOS_II_data_master_waitrequest                 (nios_ii_data_master_waitrequest),                                   //                                    .waitrequest
		.NIOS_II_data_master_byteenable                  (nios_ii_data_master_byteenable),                                    //                                    .byteenable
		.NIOS_II_data_master_read                        (nios_ii_data_master_read),                                          //                                    .read
		.NIOS_II_data_master_readdata                    (nios_ii_data_master_readdata),                                      //                                    .readdata
		.NIOS_II_data_master_write                       (nios_ii_data_master_write),                                         //                                    .write
		.NIOS_II_data_master_writedata                   (nios_ii_data_master_writedata),                                     //                                    .writedata
		.NIOS_II_data_master_debugaccess                 (nios_ii_data_master_debugaccess),                                   //                                    .debugaccess
		.NIOS_II_instruction_master_address              (nios_ii_instruction_master_address),                                //          NIOS_II_instruction_master.address
		.NIOS_II_instruction_master_waitrequest          (nios_ii_instruction_master_waitrequest),                            //                                    .waitrequest
		.NIOS_II_instruction_master_read                 (nios_ii_instruction_master_read),                                   //                                    .read
		.NIOS_II_instruction_master_readdata             (nios_ii_instruction_master_readdata),                               //                                    .readdata
		.JTAG_UART_avalon_jtag_slave_address             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),             //         JTAG_UART_avalon_jtag_slave.address
		.JTAG_UART_avalon_jtag_slave_write               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),               //                                    .write
		.JTAG_UART_avalon_jtag_slave_read                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                //                                    .read
		.JTAG_UART_avalon_jtag_slave_readdata            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),            //                                    .readdata
		.JTAG_UART_avalon_jtag_slave_writedata           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),           //                                    .writedata
		.JTAG_UART_avalon_jtag_slave_waitrequest         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),         //                                    .waitrequest
		.JTAG_UART_avalon_jtag_slave_chipselect          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),          //                                    .chipselect
		.NIOS_II_debug_mem_slave_address                 (mm_interconnect_0_nios_ii_debug_mem_slave_address),                 //             NIOS_II_debug_mem_slave.address
		.NIOS_II_debug_mem_slave_write                   (mm_interconnect_0_nios_ii_debug_mem_slave_write),                   //                                    .write
		.NIOS_II_debug_mem_slave_read                    (mm_interconnect_0_nios_ii_debug_mem_slave_read),                    //                                    .read
		.NIOS_II_debug_mem_slave_readdata                (mm_interconnect_0_nios_ii_debug_mem_slave_readdata),                //                                    .readdata
		.NIOS_II_debug_mem_slave_writedata               (mm_interconnect_0_nios_ii_debug_mem_slave_writedata),               //                                    .writedata
		.NIOS_II_debug_mem_slave_byteenable              (mm_interconnect_0_nios_ii_debug_mem_slave_byteenable),              //                                    .byteenable
		.NIOS_II_debug_mem_slave_waitrequest             (mm_interconnect_0_nios_ii_debug_mem_slave_waitrequest),             //                                    .waitrequest
		.NIOS_II_debug_mem_slave_debugaccess             (mm_interconnect_0_nios_ii_debug_mem_slave_debugaccess),             //                                    .debugaccess
		.PERFORMANCE_COUNTER_control_slave_address       (mm_interconnect_0_performance_counter_control_slave_address),       //   PERFORMANCE_COUNTER_control_slave.address
		.PERFORMANCE_COUNTER_control_slave_write         (mm_interconnect_0_performance_counter_control_slave_write),         //                                    .write
		.PERFORMANCE_COUNTER_control_slave_readdata      (mm_interconnect_0_performance_counter_control_slave_readdata),      //                                    .readdata
		.PERFORMANCE_COUNTER_control_slave_writedata     (mm_interconnect_0_performance_counter_control_slave_writedata),     //                                    .writedata
		.PERFORMANCE_COUNTER_control_slave_begintransfer (mm_interconnect_0_performance_counter_control_slave_begintransfer), //                                    .begintransfer
		.RAM_s1_address                                  (mm_interconnect_0_ram_s1_address),                                  //                              RAM_s1.address
		.RAM_s1_write                                    (mm_interconnect_0_ram_s1_write),                                    //                                    .write
		.RAM_s1_readdata                                 (mm_interconnect_0_ram_s1_readdata),                                 //                                    .readdata
		.RAM_s1_writedata                                (mm_interconnect_0_ram_s1_writedata),                                //                                    .writedata
		.RAM_s1_byteenable                               (mm_interconnect_0_ram_s1_byteenable),                               //                                    .byteenable
		.RAM_s1_chipselect                               (mm_interconnect_0_ram_s1_chipselect),                               //                                    .chipselect
		.RAM_s1_clken                                    (mm_interconnect_0_ram_s1_clken)                                     //                                    .clken
	);

	Nios2_accelerator_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios_ii_irq_irq)                 //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (nios_ii_debug_reset_request_reset),  // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
